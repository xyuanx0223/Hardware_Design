class transaction;
randc bit [3:0] a;
randc bit [3:0] b;
endclass
 
class generator;
transaction t;
mailbox mbx;
event done;
integer i;
 
function new(mailbox mbx);
this.mbx = mbx;
endfunction
 
task main();
for(i = 0; i <10; i++)begin
t = new();
t.randomize();
mbx.put(t);
$display("[GEN] :  Send Data to Driver");
  $display("SEND data: %0d & %0d", t.a, t.b);
#1;
end
->done;
endtask
endclass
 
class driver;
mailbox mbx;
transaction t;
 
function new(mailbox mbx);
this.mbx = mbx;
endfunction
 
task main();
forever begin
t = new();
mbx.get(t);
$display("[DRV] : Rcvd Data from Generator");
$display("RCVD data: %0d & %0d", t.a, t.b);
#1;
end
endtask
endclass
 
module tb();
 
transaction t;
generator gen;
driver drv;
mailbox mbx;
 
initial begin
mbx = new();
gen = new(mbx);
drv = new(mbx);
$display("----------------------------");
fork
gen.main();
drv.main();
join_any
wait(gen.done.triggered);
$display("----------------------------");
$dumpfile("dump.vcd"); 
$dumpvars;
end
endmodule
